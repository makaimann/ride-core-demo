`define ORIGINAL_MODE  3'b000
`define WAIT1_MODE     3'b001
`define DUP_MODE       3'b010
`define WAIT2_MODE     3'b011
`define CHECK_MODE     3'b100
