// Copyright (c) Stanford University
//
// This source code is patent protected and being made available under the
// terms explained in the LICENSE file in this directory.

`define ORIGINAL_MODE  3'b000
`define WAIT1_MODE     3'b001
`define DUP_MODE       3'b010
`define WAIT2_MODE     3'b011
`define CHECK_MODE     3'b100
